`timescale 1ns / 1ps

module InstMem (input [5:0] addr, output [31:0] data_out);

 reg [31:0] mem [0:63];
initial begin
    ////Experiment 1
//    mem[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
//    mem[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
//    mem[2]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
//    mem[3]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
//    mem[4]=32'b0_000000_00011_00100_000_0100_0_1100011; //beq x4, x3, 4
//    mem[5]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
//    mem[6]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
//    mem[7]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
//    mem[8]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
//    mem[9]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
//    mem[10]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
//    mem[11]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
//    mem[12]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
    //////Experiment 2
    ////mem[0] = 32'b00000000000000000_0010001010000011; //lw x5, 0(x0)
    ////mem[1] = 32'b00000000001000000_0010001100000011; //lw x6, 4(x0)
    ////mem[2] = 32'b00000000010000000_0010001110000011;  //lw x7, 8(x0)
    ////mem[3] = 32'b00100000001010011_0000001100110011;   //sub x6, x6, x5
    ////mem[4] = 32'b00000000000000011_0000010001100011;  //beq x6, x0, 8
    ////mem[5] = 32'b01111111000000000_0000110011100011;  //beq  x0, x0, -8
    ////mem[6] = 32'b00000000001010011_1000001110110011;  //add x7, x7, x5
    ////mem[7] = 32'b00000000001110000_0010100000100011;  // sw x7, 16(x0)
    //-----------------------------------------------------------------
    mem[0]=32'b0000000_00000_00000_000_00000_0110011 ;  
    mem[1]=32'h00300093 ;                               
    mem[2]=32'hffc0a113 ;                               
    mem[3]=32'h0050b193 ;                               
    mem[4]=32'hffb0b213 ;                              
    mem[5]=32'hffd0c293 ;                               
    mem[6]=32'h0040e313 ;                               
    mem[7]=32'hfff0f393 ;                               
    mem[8]=32'h00609413 ;                              
    mem[9]=32'h0020d493 ;  
    mem[10]=32'hffd00093 ;                        
    mem[11]=32'h4020d513 ; ; 
 end
 
 assign data_out = mem[addr];

endmodule